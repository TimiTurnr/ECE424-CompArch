--
-- Template
--

library ieee;
use ieee.std_logic_1164.all;


ENTITY XXX IS
    PORT(    );
END XXX;


architecture YYY of XXX is
  
 signal ZZZ;
  
BEGIN
    
END YYY;